class mem_common;
  static int num_matches;
  static int mismatches; 
endclass
